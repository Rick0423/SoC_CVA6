// Copyright 2023 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Thomas Benz <paulsc@iis.ee.ethz.ch>
// Paul Scheffler <paulsc@iis.ee.ethz.ch>
// Changed by: Mingxuan Li <mingxuanli_siris@163.com> [Peking University]

module hyperbus_delay (in_i, delay_i, out_o);
    input in_i;
    input [1:0] delay_i;
    output out_o;
    wire in_i;
    wire [1:0] delay_i;
    wire out_o;
    wire [511:0] delay_chain;
    MUX4D4BWP7T30P140 delay_mux (.I0(delay_chain[63]), .I1(delay_chain[127]), .I2(delay_chain[255]), .I3(delay_chain[511]), .S0(delay_i[0]), .S1(delay_i[1]), .Z(out_o));
    BUFFD20BWP7T30P140 delay_inst0 (.I(in_i), .Z(delay_chain[0]));
    BUFFD20BWP7T30P140 delay_inst1 (.I(delay_chain[0]), .Z(delay_chain[1]));
    BUFFD20BWP7T30P140 delay_inst2 (.I(delay_chain[1]), .Z(delay_chain[2]));
    BUFFD20BWP7T30P140 delay_inst3 (.I(delay_chain[2]), .Z(delay_chain[3]));
    BUFFD20BWP7T30P140 delay_inst4 (.I(delay_chain[3]), .Z(delay_chain[4]));
    BUFFD20BWP7T30P140 delay_inst5 (.I(delay_chain[4]), .Z(delay_chain[5]));
    BUFFD20BWP7T30P140 delay_inst6 (.I(delay_chain[5]), .Z(delay_chain[6]));
    BUFFD20BWP7T30P140 delay_inst7 (.I(delay_chain[6]), .Z(delay_chain[7]));
    BUFFD20BWP7T30P140 delay_inst8 (.I(delay_chain[7]), .Z(delay_chain[8]));
    BUFFD20BWP7T30P140 delay_inst9 (.I(delay_chain[8]), .Z(delay_chain[9]));
    BUFFD20BWP7T30P140 delay_inst10 (.I(delay_chain[9]), .Z(delay_chain[10]));
    BUFFD20BWP7T30P140 delay_inst11 (.I(delay_chain[10]), .Z(delay_chain[11]));
    BUFFD20BWP7T30P140 delay_inst12 (.I(delay_chain[11]), .Z(delay_chain[12]));
    BUFFD20BWP7T30P140 delay_inst13 (.I(delay_chain[12]), .Z(delay_chain[13]));
    BUFFD20BWP7T30P140 delay_inst14 (.I(delay_chain[13]), .Z(delay_chain[14]));
    BUFFD20BWP7T30P140 delay_inst15 (.I(delay_chain[14]), .Z(delay_chain[15]));
    BUFFD20BWP7T30P140 delay_inst16 (.I(delay_chain[15]), .Z(delay_chain[16]));
    BUFFD20BWP7T30P140 delay_inst17 (.I(delay_chain[16]), .Z(delay_chain[17]));
    BUFFD20BWP7T30P140 delay_inst18 (.I(delay_chain[17]), .Z(delay_chain[18]));
    BUFFD20BWP7T30P140 delay_inst19 (.I(delay_chain[18]), .Z(delay_chain[19]));
    BUFFD20BWP7T30P140 delay_inst20 (.I(delay_chain[19]), .Z(delay_chain[20]));
    BUFFD20BWP7T30P140 delay_inst21 (.I(delay_chain[20]), .Z(delay_chain[21]));
    BUFFD20BWP7T30P140 delay_inst22 (.I(delay_chain[21]), .Z(delay_chain[22]));
    BUFFD20BWP7T30P140 delay_inst23 (.I(delay_chain[22]), .Z(delay_chain[23]));
    BUFFD20BWP7T30P140 delay_inst24 (.I(delay_chain[23]), .Z(delay_chain[24]));
    BUFFD20BWP7T30P140 delay_inst25 (.I(delay_chain[24]), .Z(delay_chain[25]));
    BUFFD20BWP7T30P140 delay_inst26 (.I(delay_chain[25]), .Z(delay_chain[26]));
    BUFFD20BWP7T30P140 delay_inst27 (.I(delay_chain[26]), .Z(delay_chain[27]));
    BUFFD20BWP7T30P140 delay_inst28 (.I(delay_chain[27]), .Z(delay_chain[28]));
    BUFFD20BWP7T30P140 delay_inst29 (.I(delay_chain[28]), .Z(delay_chain[29]));
    BUFFD20BWP7T30P140 delay_inst30 (.I(delay_chain[29]), .Z(delay_chain[30]));
    BUFFD20BWP7T30P140 delay_inst31 (.I(delay_chain[30]), .Z(delay_chain[31]));
    BUFFD20BWP7T30P140 delay_inst32 (.I(delay_chain[31]), .Z(delay_chain[32]));
    BUFFD20BWP7T30P140 delay_inst33 (.I(delay_chain[32]), .Z(delay_chain[33]));
    BUFFD20BWP7T30P140 delay_inst34 (.I(delay_chain[33]), .Z(delay_chain[34]));
    BUFFD20BWP7T30P140 delay_inst35 (.I(delay_chain[34]), .Z(delay_chain[35]));
    BUFFD20BWP7T30P140 delay_inst36 (.I(delay_chain[35]), .Z(delay_chain[36]));
    BUFFD20BWP7T30P140 delay_inst37 (.I(delay_chain[36]), .Z(delay_chain[37]));
    BUFFD20BWP7T30P140 delay_inst38 (.I(delay_chain[37]), .Z(delay_chain[38]));
    BUFFD20BWP7T30P140 delay_inst39 (.I(delay_chain[38]), .Z(delay_chain[39]));
    BUFFD20BWP7T30P140 delay_inst40 (.I(delay_chain[39]), .Z(delay_chain[40]));
    BUFFD20BWP7T30P140 delay_inst41 (.I(delay_chain[40]), .Z(delay_chain[41]));
    BUFFD20BWP7T30P140 delay_inst42 (.I(delay_chain[41]), .Z(delay_chain[42]));
    BUFFD20BWP7T30P140 delay_inst43 (.I(delay_chain[42]), .Z(delay_chain[43]));
    BUFFD20BWP7T30P140 delay_inst44 (.I(delay_chain[43]), .Z(delay_chain[44]));
    BUFFD20BWP7T30P140 delay_inst45 (.I(delay_chain[44]), .Z(delay_chain[45]));
    BUFFD20BWP7T30P140 delay_inst46 (.I(delay_chain[45]), .Z(delay_chain[46]));
    BUFFD20BWP7T30P140 delay_inst47 (.I(delay_chain[46]), .Z(delay_chain[47]));
    BUFFD20BWP7T30P140 delay_inst48 (.I(delay_chain[47]), .Z(delay_chain[48]));
    BUFFD20BWP7T30P140 delay_inst49 (.I(delay_chain[48]), .Z(delay_chain[49]));
    BUFFD20BWP7T30P140 delay_inst50 (.I(delay_chain[49]), .Z(delay_chain[50]));
    BUFFD20BWP7T30P140 delay_inst51 (.I(delay_chain[50]), .Z(delay_chain[51]));
    BUFFD20BWP7T30P140 delay_inst52 (.I(delay_chain[51]), .Z(delay_chain[52]));
    BUFFD20BWP7T30P140 delay_inst53 (.I(delay_chain[52]), .Z(delay_chain[53]));
    BUFFD20BWP7T30P140 delay_inst54 (.I(delay_chain[53]), .Z(delay_chain[54]));
    BUFFD20BWP7T30P140 delay_inst55 (.I(delay_chain[54]), .Z(delay_chain[55]));
    BUFFD20BWP7T30P140 delay_inst56 (.I(delay_chain[55]), .Z(delay_chain[56]));
    BUFFD20BWP7T30P140 delay_inst57 (.I(delay_chain[56]), .Z(delay_chain[57]));
    BUFFD20BWP7T30P140 delay_inst58 (.I(delay_chain[57]), .Z(delay_chain[58]));
    BUFFD20BWP7T30P140 delay_inst59 (.I(delay_chain[58]), .Z(delay_chain[59]));
    BUFFD20BWP7T30P140 delay_inst60 (.I(delay_chain[59]), .Z(delay_chain[60]));
    BUFFD20BWP7T30P140 delay_inst61 (.I(delay_chain[60]), .Z(delay_chain[61]));
    BUFFD20BWP7T30P140 delay_inst62 (.I(delay_chain[61]), .Z(delay_chain[62]));
    BUFFD20BWP7T30P140 delay_inst63 (.I(delay_chain[62]), .Z(delay_chain[63]));
    BUFFD20BWP7T30P140 delay_inst64 (.I(delay_chain[63]), .Z(delay_chain[64]));
    BUFFD20BWP7T30P140 delay_inst65 (.I(delay_chain[64]), .Z(delay_chain[65]));
    BUFFD20BWP7T30P140 delay_inst66 (.I(delay_chain[65]), .Z(delay_chain[66]));
    BUFFD20BWP7T30P140 delay_inst67 (.I(delay_chain[66]), .Z(delay_chain[67]));
    BUFFD20BWP7T30P140 delay_inst68 (.I(delay_chain[67]), .Z(delay_chain[68]));
    BUFFD20BWP7T30P140 delay_inst69 (.I(delay_chain[68]), .Z(delay_chain[69]));
    BUFFD20BWP7T30P140 delay_inst70 (.I(delay_chain[69]), .Z(delay_chain[70]));
    BUFFD20BWP7T30P140 delay_inst71 (.I(delay_chain[70]), .Z(delay_chain[71]));
    BUFFD20BWP7T30P140 delay_inst72 (.I(delay_chain[71]), .Z(delay_chain[72]));
    BUFFD20BWP7T30P140 delay_inst73 (.I(delay_chain[72]), .Z(delay_chain[73]));
    BUFFD20BWP7T30P140 delay_inst74 (.I(delay_chain[73]), .Z(delay_chain[74]));
    BUFFD20BWP7T30P140 delay_inst75 (.I(delay_chain[74]), .Z(delay_chain[75]));
    BUFFD20BWP7T30P140 delay_inst76 (.I(delay_chain[75]), .Z(delay_chain[76]));
    BUFFD20BWP7T30P140 delay_inst77 (.I(delay_chain[76]), .Z(delay_chain[77]));
    BUFFD20BWP7T30P140 delay_inst78 (.I(delay_chain[77]), .Z(delay_chain[78]));
    BUFFD20BWP7T30P140 delay_inst79 (.I(delay_chain[78]), .Z(delay_chain[79]));
    BUFFD20BWP7T30P140 delay_inst80 (.I(delay_chain[79]), .Z(delay_chain[80]));
    BUFFD20BWP7T30P140 delay_inst81 (.I(delay_chain[80]), .Z(delay_chain[81]));
    BUFFD20BWP7T30P140 delay_inst82 (.I(delay_chain[81]), .Z(delay_chain[82]));
    BUFFD20BWP7T30P140 delay_inst83 (.I(delay_chain[82]), .Z(delay_chain[83]));
    BUFFD20BWP7T30P140 delay_inst84 (.I(delay_chain[83]), .Z(delay_chain[84]));
    BUFFD20BWP7T30P140 delay_inst85 (.I(delay_chain[84]), .Z(delay_chain[85]));
    BUFFD20BWP7T30P140 delay_inst86 (.I(delay_chain[85]), .Z(delay_chain[86]));
    BUFFD20BWP7T30P140 delay_inst87 (.I(delay_chain[86]), .Z(delay_chain[87]));
    BUFFD20BWP7T30P140 delay_inst88 (.I(delay_chain[87]), .Z(delay_chain[88]));
    BUFFD20BWP7T30P140 delay_inst89 (.I(delay_chain[88]), .Z(delay_chain[89]));
    BUFFD20BWP7T30P140 delay_inst90 (.I(delay_chain[89]), .Z(delay_chain[90]));
    BUFFD20BWP7T30P140 delay_inst91 (.I(delay_chain[90]), .Z(delay_chain[91]));
    BUFFD20BWP7T30P140 delay_inst92 (.I(delay_chain[91]), .Z(delay_chain[92]));
    BUFFD20BWP7T30P140 delay_inst93 (.I(delay_chain[92]), .Z(delay_chain[93]));
    BUFFD20BWP7T30P140 delay_inst94 (.I(delay_chain[93]), .Z(delay_chain[94]));
    BUFFD20BWP7T30P140 delay_inst95 (.I(delay_chain[94]), .Z(delay_chain[95]));
    BUFFD20BWP7T30P140 delay_inst96 (.I(delay_chain[95]), .Z(delay_chain[96]));
    BUFFD20BWP7T30P140 delay_inst97 (.I(delay_chain[96]), .Z(delay_chain[97]));
    BUFFD20BWP7T30P140 delay_inst98 (.I(delay_chain[97]), .Z(delay_chain[98]));
    BUFFD20BWP7T30P140 delay_inst99 (.I(delay_chain[98]), .Z(delay_chain[99]));
    BUFFD20BWP7T30P140 delay_inst100 (.I(delay_chain[99]), .Z(delay_chain[100]));
    BUFFD20BWP7T30P140 delay_inst101 (.I(delay_chain[100]), .Z(delay_chain[101]));
    BUFFD20BWP7T30P140 delay_inst102 (.I(delay_chain[101]), .Z(delay_chain[102]));
    BUFFD20BWP7T30P140 delay_inst103 (.I(delay_chain[102]), .Z(delay_chain[103]));
    BUFFD20BWP7T30P140 delay_inst104 (.I(delay_chain[103]), .Z(delay_chain[104]));
    BUFFD20BWP7T30P140 delay_inst105 (.I(delay_chain[104]), .Z(delay_chain[105]));
    BUFFD20BWP7T30P140 delay_inst106 (.I(delay_chain[105]), .Z(delay_chain[106]));
    BUFFD20BWP7T30P140 delay_inst107 (.I(delay_chain[106]), .Z(delay_chain[107]));
    BUFFD20BWP7T30P140 delay_inst108 (.I(delay_chain[107]), .Z(delay_chain[108]));
    BUFFD20BWP7T30P140 delay_inst109 (.I(delay_chain[108]), .Z(delay_chain[109]));
    BUFFD20BWP7T30P140 delay_inst110 (.I(delay_chain[109]), .Z(delay_chain[110]));
    BUFFD20BWP7T30P140 delay_inst111 (.I(delay_chain[110]), .Z(delay_chain[111]));
    BUFFD20BWP7T30P140 delay_inst112 (.I(delay_chain[111]), .Z(delay_chain[112]));
    BUFFD20BWP7T30P140 delay_inst113 (.I(delay_chain[112]), .Z(delay_chain[113]));
    BUFFD20BWP7T30P140 delay_inst114 (.I(delay_chain[113]), .Z(delay_chain[114]));
    BUFFD20BWP7T30P140 delay_inst115 (.I(delay_chain[114]), .Z(delay_chain[115]));
    BUFFD20BWP7T30P140 delay_inst116 (.I(delay_chain[115]), .Z(delay_chain[116]));
    BUFFD20BWP7T30P140 delay_inst117 (.I(delay_chain[116]), .Z(delay_chain[117]));
    BUFFD20BWP7T30P140 delay_inst118 (.I(delay_chain[117]), .Z(delay_chain[118]));
    BUFFD20BWP7T30P140 delay_inst119 (.I(delay_chain[118]), .Z(delay_chain[119]));
    BUFFD20BWP7T30P140 delay_inst120 (.I(delay_chain[119]), .Z(delay_chain[120]));
    BUFFD20BWP7T30P140 delay_inst121 (.I(delay_chain[120]), .Z(delay_chain[121]));
    BUFFD20BWP7T30P140 delay_inst122 (.I(delay_chain[121]), .Z(delay_chain[122]));
    BUFFD20BWP7T30P140 delay_inst123 (.I(delay_chain[122]), .Z(delay_chain[123]));
    BUFFD20BWP7T30P140 delay_inst124 (.I(delay_chain[123]), .Z(delay_chain[124]));
    BUFFD20BWP7T30P140 delay_inst125 (.I(delay_chain[124]), .Z(delay_chain[125]));
    BUFFD20BWP7T30P140 delay_inst126 (.I(delay_chain[125]), .Z(delay_chain[126]));
    BUFFD20BWP7T30P140 delay_inst127 (.I(delay_chain[126]), .Z(delay_chain[127]));
    BUFFD20BWP7T30P140 delay_inst128 (.I(delay_chain[127]), .Z(delay_chain[128]));
    BUFFD20BWP7T30P140 delay_inst129 (.I(delay_chain[128]), .Z(delay_chain[129]));
    BUFFD20BWP7T30P140 delay_inst130 (.I(delay_chain[129]), .Z(delay_chain[130]));
    BUFFD20BWP7T30P140 delay_inst131 (.I(delay_chain[130]), .Z(delay_chain[131]));
    BUFFD20BWP7T30P140 delay_inst132 (.I(delay_chain[131]), .Z(delay_chain[132]));
    BUFFD20BWP7T30P140 delay_inst133 (.I(delay_chain[132]), .Z(delay_chain[133]));
    BUFFD20BWP7T30P140 delay_inst134 (.I(delay_chain[133]), .Z(delay_chain[134]));
    BUFFD20BWP7T30P140 delay_inst135 (.I(delay_chain[134]), .Z(delay_chain[135]));
    BUFFD20BWP7T30P140 delay_inst136 (.I(delay_chain[135]), .Z(delay_chain[136]));
    BUFFD20BWP7T30P140 delay_inst137 (.I(delay_chain[136]), .Z(delay_chain[137]));
    BUFFD20BWP7T30P140 delay_inst138 (.I(delay_chain[137]), .Z(delay_chain[138]));
    BUFFD20BWP7T30P140 delay_inst139 (.I(delay_chain[138]), .Z(delay_chain[139]));
    BUFFD20BWP7T30P140 delay_inst140 (.I(delay_chain[139]), .Z(delay_chain[140]));
    BUFFD20BWP7T30P140 delay_inst141 (.I(delay_chain[140]), .Z(delay_chain[141]));
    BUFFD20BWP7T30P140 delay_inst142 (.I(delay_chain[141]), .Z(delay_chain[142]));
    BUFFD20BWP7T30P140 delay_inst143 (.I(delay_chain[142]), .Z(delay_chain[143]));
    BUFFD20BWP7T30P140 delay_inst144 (.I(delay_chain[143]), .Z(delay_chain[144]));
    BUFFD20BWP7T30P140 delay_inst145 (.I(delay_chain[144]), .Z(delay_chain[145]));
    BUFFD20BWP7T30P140 delay_inst146 (.I(delay_chain[145]), .Z(delay_chain[146]));
    BUFFD20BWP7T30P140 delay_inst147 (.I(delay_chain[146]), .Z(delay_chain[147]));
    BUFFD20BWP7T30P140 delay_inst148 (.I(delay_chain[147]), .Z(delay_chain[148]));
    BUFFD20BWP7T30P140 delay_inst149 (.I(delay_chain[148]), .Z(delay_chain[149]));
    BUFFD20BWP7T30P140 delay_inst150 (.I(delay_chain[149]), .Z(delay_chain[150]));
    BUFFD20BWP7T30P140 delay_inst151 (.I(delay_chain[150]), .Z(delay_chain[151]));
    BUFFD20BWP7T30P140 delay_inst152 (.I(delay_chain[151]), .Z(delay_chain[152]));
    BUFFD20BWP7T30P140 delay_inst153 (.I(delay_chain[152]), .Z(delay_chain[153]));
    BUFFD20BWP7T30P140 delay_inst154 (.I(delay_chain[153]), .Z(delay_chain[154]));
    BUFFD20BWP7T30P140 delay_inst155 (.I(delay_chain[154]), .Z(delay_chain[155]));
    BUFFD20BWP7T30P140 delay_inst156 (.I(delay_chain[155]), .Z(delay_chain[156]));
    BUFFD20BWP7T30P140 delay_inst157 (.I(delay_chain[156]), .Z(delay_chain[157]));
    BUFFD20BWP7T30P140 delay_inst158 (.I(delay_chain[157]), .Z(delay_chain[158]));
    BUFFD20BWP7T30P140 delay_inst159 (.I(delay_chain[158]), .Z(delay_chain[159]));
    BUFFD20BWP7T30P140 delay_inst160 (.I(delay_chain[159]), .Z(delay_chain[160]));
    BUFFD20BWP7T30P140 delay_inst161 (.I(delay_chain[160]), .Z(delay_chain[161]));
    BUFFD20BWP7T30P140 delay_inst162 (.I(delay_chain[161]), .Z(delay_chain[162]));
    BUFFD20BWP7T30P140 delay_inst163 (.I(delay_chain[162]), .Z(delay_chain[163]));
    BUFFD20BWP7T30P140 delay_inst164 (.I(delay_chain[163]), .Z(delay_chain[164]));
    BUFFD20BWP7T30P140 delay_inst165 (.I(delay_chain[164]), .Z(delay_chain[165]));
    BUFFD20BWP7T30P140 delay_inst166 (.I(delay_chain[165]), .Z(delay_chain[166]));
    BUFFD20BWP7T30P140 delay_inst167 (.I(delay_chain[166]), .Z(delay_chain[167]));
    BUFFD20BWP7T30P140 delay_inst168 (.I(delay_chain[167]), .Z(delay_chain[168]));
    BUFFD20BWP7T30P140 delay_inst169 (.I(delay_chain[168]), .Z(delay_chain[169]));
    BUFFD20BWP7T30P140 delay_inst170 (.I(delay_chain[169]), .Z(delay_chain[170]));
    BUFFD20BWP7T30P140 delay_inst171 (.I(delay_chain[170]), .Z(delay_chain[171]));
    BUFFD20BWP7T30P140 delay_inst172 (.I(delay_chain[171]), .Z(delay_chain[172]));
    BUFFD20BWP7T30P140 delay_inst173 (.I(delay_chain[172]), .Z(delay_chain[173]));
    BUFFD20BWP7T30P140 delay_inst174 (.I(delay_chain[173]), .Z(delay_chain[174]));
    BUFFD20BWP7T30P140 delay_inst175 (.I(delay_chain[174]), .Z(delay_chain[175]));
    BUFFD20BWP7T30P140 delay_inst176 (.I(delay_chain[175]), .Z(delay_chain[176]));
    BUFFD20BWP7T30P140 delay_inst177 (.I(delay_chain[176]), .Z(delay_chain[177]));
    BUFFD20BWP7T30P140 delay_inst178 (.I(delay_chain[177]), .Z(delay_chain[178]));
    BUFFD20BWP7T30P140 delay_inst179 (.I(delay_chain[178]), .Z(delay_chain[179]));
    BUFFD20BWP7T30P140 delay_inst180 (.I(delay_chain[179]), .Z(delay_chain[180]));
    BUFFD20BWP7T30P140 delay_inst181 (.I(delay_chain[180]), .Z(delay_chain[181]));
    BUFFD20BWP7T30P140 delay_inst182 (.I(delay_chain[181]), .Z(delay_chain[182]));
    BUFFD20BWP7T30P140 delay_inst183 (.I(delay_chain[182]), .Z(delay_chain[183]));
    BUFFD20BWP7T30P140 delay_inst184 (.I(delay_chain[183]), .Z(delay_chain[184]));
    BUFFD20BWP7T30P140 delay_inst185 (.I(delay_chain[184]), .Z(delay_chain[185]));
    BUFFD20BWP7T30P140 delay_inst186 (.I(delay_chain[185]), .Z(delay_chain[186]));
    BUFFD20BWP7T30P140 delay_inst187 (.I(delay_chain[186]), .Z(delay_chain[187]));
    BUFFD20BWP7T30P140 delay_inst188 (.I(delay_chain[187]), .Z(delay_chain[188]));
    BUFFD20BWP7T30P140 delay_inst189 (.I(delay_chain[188]), .Z(delay_chain[189]));
    BUFFD20BWP7T30P140 delay_inst190 (.I(delay_chain[189]), .Z(delay_chain[190]));
    BUFFD20BWP7T30P140 delay_inst191 (.I(delay_chain[190]), .Z(delay_chain[191]));
    BUFFD20BWP7T30P140 delay_inst192 (.I(delay_chain[191]), .Z(delay_chain[192]));
    BUFFD20BWP7T30P140 delay_inst193 (.I(delay_chain[192]), .Z(delay_chain[193]));
    BUFFD20BWP7T30P140 delay_inst194 (.I(delay_chain[193]), .Z(delay_chain[194]));
    BUFFD20BWP7T30P140 delay_inst195 (.I(delay_chain[194]), .Z(delay_chain[195]));
    BUFFD20BWP7T30P140 delay_inst196 (.I(delay_chain[195]), .Z(delay_chain[196]));
    BUFFD20BWP7T30P140 delay_inst197 (.I(delay_chain[196]), .Z(delay_chain[197]));
    BUFFD20BWP7T30P140 delay_inst198 (.I(delay_chain[197]), .Z(delay_chain[198]));
    BUFFD20BWP7T30P140 delay_inst199 (.I(delay_chain[198]), .Z(delay_chain[199]));
    BUFFD20BWP7T30P140 delay_inst200 (.I(delay_chain[199]), .Z(delay_chain[200]));
    BUFFD20BWP7T30P140 delay_inst201 (.I(delay_chain[200]), .Z(delay_chain[201]));
    BUFFD20BWP7T30P140 delay_inst202 (.I(delay_chain[201]), .Z(delay_chain[202]));
    BUFFD20BWP7T30P140 delay_inst203 (.I(delay_chain[202]), .Z(delay_chain[203]));
    BUFFD20BWP7T30P140 delay_inst204 (.I(delay_chain[203]), .Z(delay_chain[204]));
    BUFFD20BWP7T30P140 delay_inst205 (.I(delay_chain[204]), .Z(delay_chain[205]));
    BUFFD20BWP7T30P140 delay_inst206 (.I(delay_chain[205]), .Z(delay_chain[206]));
    BUFFD20BWP7T30P140 delay_inst207 (.I(delay_chain[206]), .Z(delay_chain[207]));
    BUFFD20BWP7T30P140 delay_inst208 (.I(delay_chain[207]), .Z(delay_chain[208]));
    BUFFD20BWP7T30P140 delay_inst209 (.I(delay_chain[208]), .Z(delay_chain[209]));
    BUFFD20BWP7T30P140 delay_inst210 (.I(delay_chain[209]), .Z(delay_chain[210]));
    BUFFD20BWP7T30P140 delay_inst211 (.I(delay_chain[210]), .Z(delay_chain[211]));
    BUFFD20BWP7T30P140 delay_inst212 (.I(delay_chain[211]), .Z(delay_chain[212]));
    BUFFD20BWP7T30P140 delay_inst213 (.I(delay_chain[212]), .Z(delay_chain[213]));
    BUFFD20BWP7T30P140 delay_inst214 (.I(delay_chain[213]), .Z(delay_chain[214]));
    BUFFD20BWP7T30P140 delay_inst215 (.I(delay_chain[214]), .Z(delay_chain[215]));
    BUFFD20BWP7T30P140 delay_inst216 (.I(delay_chain[215]), .Z(delay_chain[216]));
    BUFFD20BWP7T30P140 delay_inst217 (.I(delay_chain[216]), .Z(delay_chain[217]));
    BUFFD20BWP7T30P140 delay_inst218 (.I(delay_chain[217]), .Z(delay_chain[218]));
    BUFFD20BWP7T30P140 delay_inst219 (.I(delay_chain[218]), .Z(delay_chain[219]));
    BUFFD20BWP7T30P140 delay_inst220 (.I(delay_chain[219]), .Z(delay_chain[220]));
    BUFFD20BWP7T30P140 delay_inst221 (.I(delay_chain[220]), .Z(delay_chain[221]));
    BUFFD20BWP7T30P140 delay_inst222 (.I(delay_chain[221]), .Z(delay_chain[222]));
    BUFFD20BWP7T30P140 delay_inst223 (.I(delay_chain[222]), .Z(delay_chain[223]));
    BUFFD20BWP7T30P140 delay_inst224 (.I(delay_chain[223]), .Z(delay_chain[224]));
    BUFFD20BWP7T30P140 delay_inst225 (.I(delay_chain[224]), .Z(delay_chain[225]));
    BUFFD20BWP7T30P140 delay_inst226 (.I(delay_chain[225]), .Z(delay_chain[226]));
    BUFFD20BWP7T30P140 delay_inst227 (.I(delay_chain[226]), .Z(delay_chain[227]));
    BUFFD20BWP7T30P140 delay_inst228 (.I(delay_chain[227]), .Z(delay_chain[228]));
    BUFFD20BWP7T30P140 delay_inst229 (.I(delay_chain[228]), .Z(delay_chain[229]));
    BUFFD20BWP7T30P140 delay_inst230 (.I(delay_chain[229]), .Z(delay_chain[230]));
    BUFFD20BWP7T30P140 delay_inst231 (.I(delay_chain[230]), .Z(delay_chain[231]));
    BUFFD20BWP7T30P140 delay_inst232 (.I(delay_chain[231]), .Z(delay_chain[232]));
    BUFFD20BWP7T30P140 delay_inst233 (.I(delay_chain[232]), .Z(delay_chain[233]));
    BUFFD20BWP7T30P140 delay_inst234 (.I(delay_chain[233]), .Z(delay_chain[234]));
    BUFFD20BWP7T30P140 delay_inst235 (.I(delay_chain[234]), .Z(delay_chain[235]));
    BUFFD20BWP7T30P140 delay_inst236 (.I(delay_chain[235]), .Z(delay_chain[236]));
    BUFFD20BWP7T30P140 delay_inst237 (.I(delay_chain[236]), .Z(delay_chain[237]));
    BUFFD20BWP7T30P140 delay_inst238 (.I(delay_chain[237]), .Z(delay_chain[238]));
    BUFFD20BWP7T30P140 delay_inst239 (.I(delay_chain[238]), .Z(delay_chain[239]));
    BUFFD20BWP7T30P140 delay_inst240 (.I(delay_chain[239]), .Z(delay_chain[240]));
    BUFFD20BWP7T30P140 delay_inst241 (.I(delay_chain[240]), .Z(delay_chain[241]));
    BUFFD20BWP7T30P140 delay_inst242 (.I(delay_chain[241]), .Z(delay_chain[242]));
    BUFFD20BWP7T30P140 delay_inst243 (.I(delay_chain[242]), .Z(delay_chain[243]));
    BUFFD20BWP7T30P140 delay_inst244 (.I(delay_chain[243]), .Z(delay_chain[244]));
    BUFFD20BWP7T30P140 delay_inst245 (.I(delay_chain[244]), .Z(delay_chain[245]));
    BUFFD20BWP7T30P140 delay_inst246 (.I(delay_chain[245]), .Z(delay_chain[246]));
    BUFFD20BWP7T30P140 delay_inst247 (.I(delay_chain[246]), .Z(delay_chain[247]));
    BUFFD20BWP7T30P140 delay_inst248 (.I(delay_chain[247]), .Z(delay_chain[248]));
    BUFFD20BWP7T30P140 delay_inst249 (.I(delay_chain[248]), .Z(delay_chain[249]));
    BUFFD20BWP7T30P140 delay_inst250 (.I(delay_chain[249]), .Z(delay_chain[250]));
    BUFFD20BWP7T30P140 delay_inst251 (.I(delay_chain[250]), .Z(delay_chain[251]));
    BUFFD20BWP7T30P140 delay_inst252 (.I(delay_chain[251]), .Z(delay_chain[252]));
    BUFFD20BWP7T30P140 delay_inst253 (.I(delay_chain[252]), .Z(delay_chain[253]));
    BUFFD20BWP7T30P140 delay_inst254 (.I(delay_chain[253]), .Z(delay_chain[254]));
    BUFFD20BWP7T30P140 delay_inst255 (.I(delay_chain[254]), .Z(delay_chain[255]));
    BUFFD20BWP7T30P140 delay_inst256 (.I(delay_chain[255]), .Z(delay_chain[256]));
    BUFFD20BWP7T30P140 delay_inst257 (.I(delay_chain[256]), .Z(delay_chain[257]));
    BUFFD20BWP7T30P140 delay_inst258 (.I(delay_chain[257]), .Z(delay_chain[258]));
    BUFFD20BWP7T30P140 delay_inst259 (.I(delay_chain[258]), .Z(delay_chain[259]));
    BUFFD20BWP7T30P140 delay_inst260 (.I(delay_chain[259]), .Z(delay_chain[260]));
    BUFFD20BWP7T30P140 delay_inst261 (.I(delay_chain[260]), .Z(delay_chain[261]));
    BUFFD20BWP7T30P140 delay_inst262 (.I(delay_chain[261]), .Z(delay_chain[262]));
    BUFFD20BWP7T30P140 delay_inst263 (.I(delay_chain[262]), .Z(delay_chain[263]));
    BUFFD20BWP7T30P140 delay_inst264 (.I(delay_chain[263]), .Z(delay_chain[264]));
    BUFFD20BWP7T30P140 delay_inst265 (.I(delay_chain[264]), .Z(delay_chain[265]));
    BUFFD20BWP7T30P140 delay_inst266 (.I(delay_chain[265]), .Z(delay_chain[266]));
    BUFFD20BWP7T30P140 delay_inst267 (.I(delay_chain[266]), .Z(delay_chain[267]));
    BUFFD20BWP7T30P140 delay_inst268 (.I(delay_chain[267]), .Z(delay_chain[268]));
    BUFFD20BWP7T30P140 delay_inst269 (.I(delay_chain[268]), .Z(delay_chain[269]));
    BUFFD20BWP7T30P140 delay_inst270 (.I(delay_chain[269]), .Z(delay_chain[270]));
    BUFFD20BWP7T30P140 delay_inst271 (.I(delay_chain[270]), .Z(delay_chain[271]));
    BUFFD20BWP7T30P140 delay_inst272 (.I(delay_chain[271]), .Z(delay_chain[272]));
    BUFFD20BWP7T30P140 delay_inst273 (.I(delay_chain[272]), .Z(delay_chain[273]));
    BUFFD20BWP7T30P140 delay_inst274 (.I(delay_chain[273]), .Z(delay_chain[274]));
    BUFFD20BWP7T30P140 delay_inst275 (.I(delay_chain[274]), .Z(delay_chain[275]));
    BUFFD20BWP7T30P140 delay_inst276 (.I(delay_chain[275]), .Z(delay_chain[276]));
    BUFFD20BWP7T30P140 delay_inst277 (.I(delay_chain[276]), .Z(delay_chain[277]));
    BUFFD20BWP7T30P140 delay_inst278 (.I(delay_chain[277]), .Z(delay_chain[278]));
    BUFFD20BWP7T30P140 delay_inst279 (.I(delay_chain[278]), .Z(delay_chain[279]));
    BUFFD20BWP7T30P140 delay_inst280 (.I(delay_chain[279]), .Z(delay_chain[280]));
    BUFFD20BWP7T30P140 delay_inst281 (.I(delay_chain[280]), .Z(delay_chain[281]));
    BUFFD20BWP7T30P140 delay_inst282 (.I(delay_chain[281]), .Z(delay_chain[282]));
    BUFFD20BWP7T30P140 delay_inst283 (.I(delay_chain[282]), .Z(delay_chain[283]));
    BUFFD20BWP7T30P140 delay_inst284 (.I(delay_chain[283]), .Z(delay_chain[284]));
    BUFFD20BWP7T30P140 delay_inst285 (.I(delay_chain[284]), .Z(delay_chain[285]));
    BUFFD20BWP7T30P140 delay_inst286 (.I(delay_chain[285]), .Z(delay_chain[286]));
    BUFFD20BWP7T30P140 delay_inst287 (.I(delay_chain[286]), .Z(delay_chain[287]));
    BUFFD20BWP7T30P140 delay_inst288 (.I(delay_chain[287]), .Z(delay_chain[288]));
    BUFFD20BWP7T30P140 delay_inst289 (.I(delay_chain[288]), .Z(delay_chain[289]));
    BUFFD20BWP7T30P140 delay_inst290 (.I(delay_chain[289]), .Z(delay_chain[290]));
    BUFFD20BWP7T30P140 delay_inst291 (.I(delay_chain[290]), .Z(delay_chain[291]));
    BUFFD20BWP7T30P140 delay_inst292 (.I(delay_chain[291]), .Z(delay_chain[292]));
    BUFFD20BWP7T30P140 delay_inst293 (.I(delay_chain[292]), .Z(delay_chain[293]));
    BUFFD20BWP7T30P140 delay_inst294 (.I(delay_chain[293]), .Z(delay_chain[294]));
    BUFFD20BWP7T30P140 delay_inst295 (.I(delay_chain[294]), .Z(delay_chain[295]));
    BUFFD20BWP7T30P140 delay_inst296 (.I(delay_chain[295]), .Z(delay_chain[296]));
    BUFFD20BWP7T30P140 delay_inst297 (.I(delay_chain[296]), .Z(delay_chain[297]));
    BUFFD20BWP7T30P140 delay_inst298 (.I(delay_chain[297]), .Z(delay_chain[298]));
    BUFFD20BWP7T30P140 delay_inst299 (.I(delay_chain[298]), .Z(delay_chain[299]));
    BUFFD20BWP7T30P140 delay_inst300 (.I(delay_chain[299]), .Z(delay_chain[300]));
    BUFFD20BWP7T30P140 delay_inst301 (.I(delay_chain[300]), .Z(delay_chain[301]));
    BUFFD20BWP7T30P140 delay_inst302 (.I(delay_chain[301]), .Z(delay_chain[302]));
    BUFFD20BWP7T30P140 delay_inst303 (.I(delay_chain[302]), .Z(delay_chain[303]));
    BUFFD20BWP7T30P140 delay_inst304 (.I(delay_chain[303]), .Z(delay_chain[304]));
    BUFFD20BWP7T30P140 delay_inst305 (.I(delay_chain[304]), .Z(delay_chain[305]));
    BUFFD20BWP7T30P140 delay_inst306 (.I(delay_chain[305]), .Z(delay_chain[306]));
    BUFFD20BWP7T30P140 delay_inst307 (.I(delay_chain[306]), .Z(delay_chain[307]));
    BUFFD20BWP7T30P140 delay_inst308 (.I(delay_chain[307]), .Z(delay_chain[308]));
    BUFFD20BWP7T30P140 delay_inst309 (.I(delay_chain[308]), .Z(delay_chain[309]));
    BUFFD20BWP7T30P140 delay_inst310 (.I(delay_chain[309]), .Z(delay_chain[310]));
    BUFFD20BWP7T30P140 delay_inst311 (.I(delay_chain[310]), .Z(delay_chain[311]));
    BUFFD20BWP7T30P140 delay_inst312 (.I(delay_chain[311]), .Z(delay_chain[312]));
    BUFFD20BWP7T30P140 delay_inst313 (.I(delay_chain[312]), .Z(delay_chain[313]));
    BUFFD20BWP7T30P140 delay_inst314 (.I(delay_chain[313]), .Z(delay_chain[314]));
    BUFFD20BWP7T30P140 delay_inst315 (.I(delay_chain[314]), .Z(delay_chain[315]));
    BUFFD20BWP7T30P140 delay_inst316 (.I(delay_chain[315]), .Z(delay_chain[316]));
    BUFFD20BWP7T30P140 delay_inst317 (.I(delay_chain[316]), .Z(delay_chain[317]));
    BUFFD20BWP7T30P140 delay_inst318 (.I(delay_chain[317]), .Z(delay_chain[318]));
    BUFFD20BWP7T30P140 delay_inst319 (.I(delay_chain[318]), .Z(delay_chain[319]));
    BUFFD20BWP7T30P140 delay_inst320 (.I(delay_chain[319]), .Z(delay_chain[320]));
    BUFFD20BWP7T30P140 delay_inst321 (.I(delay_chain[320]), .Z(delay_chain[321]));
    BUFFD20BWP7T30P140 delay_inst322 (.I(delay_chain[321]), .Z(delay_chain[322]));
    BUFFD20BWP7T30P140 delay_inst323 (.I(delay_chain[322]), .Z(delay_chain[323]));
    BUFFD20BWP7T30P140 delay_inst324 (.I(delay_chain[323]), .Z(delay_chain[324]));
    BUFFD20BWP7T30P140 delay_inst325 (.I(delay_chain[324]), .Z(delay_chain[325]));
    BUFFD20BWP7T30P140 delay_inst326 (.I(delay_chain[325]), .Z(delay_chain[326]));
    BUFFD20BWP7T30P140 delay_inst327 (.I(delay_chain[326]), .Z(delay_chain[327]));
    BUFFD20BWP7T30P140 delay_inst328 (.I(delay_chain[327]), .Z(delay_chain[328]));
    BUFFD20BWP7T30P140 delay_inst329 (.I(delay_chain[328]), .Z(delay_chain[329]));
    BUFFD20BWP7T30P140 delay_inst330 (.I(delay_chain[329]), .Z(delay_chain[330]));
    BUFFD20BWP7T30P140 delay_inst331 (.I(delay_chain[330]), .Z(delay_chain[331]));
    BUFFD20BWP7T30P140 delay_inst332 (.I(delay_chain[331]), .Z(delay_chain[332]));
    BUFFD20BWP7T30P140 delay_inst333 (.I(delay_chain[332]), .Z(delay_chain[333]));
    BUFFD20BWP7T30P140 delay_inst334 (.I(delay_chain[333]), .Z(delay_chain[334]));
    BUFFD20BWP7T30P140 delay_inst335 (.I(delay_chain[334]), .Z(delay_chain[335]));
    BUFFD20BWP7T30P140 delay_inst336 (.I(delay_chain[335]), .Z(delay_chain[336]));
    BUFFD20BWP7T30P140 delay_inst337 (.I(delay_chain[336]), .Z(delay_chain[337]));
    BUFFD20BWP7T30P140 delay_inst338 (.I(delay_chain[337]), .Z(delay_chain[338]));
    BUFFD20BWP7T30P140 delay_inst339 (.I(delay_chain[338]), .Z(delay_chain[339]));
    BUFFD20BWP7T30P140 delay_inst340 (.I(delay_chain[339]), .Z(delay_chain[340]));
    BUFFD20BWP7T30P140 delay_inst341 (.I(delay_chain[340]), .Z(delay_chain[341]));
    BUFFD20BWP7T30P140 delay_inst342 (.I(delay_chain[341]), .Z(delay_chain[342]));
    BUFFD20BWP7T30P140 delay_inst343 (.I(delay_chain[342]), .Z(delay_chain[343]));
    BUFFD20BWP7T30P140 delay_inst344 (.I(delay_chain[343]), .Z(delay_chain[344]));
    BUFFD20BWP7T30P140 delay_inst345 (.I(delay_chain[344]), .Z(delay_chain[345]));
    BUFFD20BWP7T30P140 delay_inst346 (.I(delay_chain[345]), .Z(delay_chain[346]));
    BUFFD20BWP7T30P140 delay_inst347 (.I(delay_chain[346]), .Z(delay_chain[347]));
    BUFFD20BWP7T30P140 delay_inst348 (.I(delay_chain[347]), .Z(delay_chain[348]));
    BUFFD20BWP7T30P140 delay_inst349 (.I(delay_chain[348]), .Z(delay_chain[349]));
    BUFFD20BWP7T30P140 delay_inst350 (.I(delay_chain[349]), .Z(delay_chain[350]));
    BUFFD20BWP7T30P140 delay_inst351 (.I(delay_chain[350]), .Z(delay_chain[351]));
    BUFFD20BWP7T30P140 delay_inst352 (.I(delay_chain[351]), .Z(delay_chain[352]));
    BUFFD20BWP7T30P140 delay_inst353 (.I(delay_chain[352]), .Z(delay_chain[353]));
    BUFFD20BWP7T30P140 delay_inst354 (.I(delay_chain[353]), .Z(delay_chain[354]));
    BUFFD20BWP7T30P140 delay_inst355 (.I(delay_chain[354]), .Z(delay_chain[355]));
    BUFFD20BWP7T30P140 delay_inst356 (.I(delay_chain[355]), .Z(delay_chain[356]));
    BUFFD20BWP7T30P140 delay_inst357 (.I(delay_chain[356]), .Z(delay_chain[357]));
    BUFFD20BWP7T30P140 delay_inst358 (.I(delay_chain[357]), .Z(delay_chain[358]));
    BUFFD20BWP7T30P140 delay_inst359 (.I(delay_chain[358]), .Z(delay_chain[359]));
    BUFFD20BWP7T30P140 delay_inst360 (.I(delay_chain[359]), .Z(delay_chain[360]));
    BUFFD20BWP7T30P140 delay_inst361 (.I(delay_chain[360]), .Z(delay_chain[361]));
    BUFFD20BWP7T30P140 delay_inst362 (.I(delay_chain[361]), .Z(delay_chain[362]));
    BUFFD20BWP7T30P140 delay_inst363 (.I(delay_chain[362]), .Z(delay_chain[363]));
    BUFFD20BWP7T30P140 delay_inst364 (.I(delay_chain[363]), .Z(delay_chain[364]));
    BUFFD20BWP7T30P140 delay_inst365 (.I(delay_chain[364]), .Z(delay_chain[365]));
    BUFFD20BWP7T30P140 delay_inst366 (.I(delay_chain[365]), .Z(delay_chain[366]));
    BUFFD20BWP7T30P140 delay_inst367 (.I(delay_chain[366]), .Z(delay_chain[367]));
    BUFFD20BWP7T30P140 delay_inst368 (.I(delay_chain[367]), .Z(delay_chain[368]));
    BUFFD20BWP7T30P140 delay_inst369 (.I(delay_chain[368]), .Z(delay_chain[369]));
    BUFFD20BWP7T30P140 delay_inst370 (.I(delay_chain[369]), .Z(delay_chain[370]));
    BUFFD20BWP7T30P140 delay_inst371 (.I(delay_chain[370]), .Z(delay_chain[371]));
    BUFFD20BWP7T30P140 delay_inst372 (.I(delay_chain[371]), .Z(delay_chain[372]));
    BUFFD20BWP7T30P140 delay_inst373 (.I(delay_chain[372]), .Z(delay_chain[373]));
    BUFFD20BWP7T30P140 delay_inst374 (.I(delay_chain[373]), .Z(delay_chain[374]));
    BUFFD20BWP7T30P140 delay_inst375 (.I(delay_chain[374]), .Z(delay_chain[375]));
    BUFFD20BWP7T30P140 delay_inst376 (.I(delay_chain[375]), .Z(delay_chain[376]));
    BUFFD20BWP7T30P140 delay_inst377 (.I(delay_chain[376]), .Z(delay_chain[377]));
    BUFFD20BWP7T30P140 delay_inst378 (.I(delay_chain[377]), .Z(delay_chain[378]));
    BUFFD20BWP7T30P140 delay_inst379 (.I(delay_chain[378]), .Z(delay_chain[379]));
    BUFFD20BWP7T30P140 delay_inst380 (.I(delay_chain[379]), .Z(delay_chain[380]));
    BUFFD20BWP7T30P140 delay_inst381 (.I(delay_chain[380]), .Z(delay_chain[381]));
    BUFFD20BWP7T30P140 delay_inst382 (.I(delay_chain[381]), .Z(delay_chain[382]));
    BUFFD20BWP7T30P140 delay_inst383 (.I(delay_chain[382]), .Z(delay_chain[383]));
    BUFFD20BWP7T30P140 delay_inst384 (.I(delay_chain[383]), .Z(delay_chain[384]));
    BUFFD20BWP7T30P140 delay_inst385 (.I(delay_chain[384]), .Z(delay_chain[385]));
    BUFFD20BWP7T30P140 delay_inst386 (.I(delay_chain[385]), .Z(delay_chain[386]));
    BUFFD20BWP7T30P140 delay_inst387 (.I(delay_chain[386]), .Z(delay_chain[387]));
    BUFFD20BWP7T30P140 delay_inst388 (.I(delay_chain[387]), .Z(delay_chain[388]));
    BUFFD20BWP7T30P140 delay_inst389 (.I(delay_chain[388]), .Z(delay_chain[389]));
    BUFFD20BWP7T30P140 delay_inst390 (.I(delay_chain[389]), .Z(delay_chain[390]));
    BUFFD20BWP7T30P140 delay_inst391 (.I(delay_chain[390]), .Z(delay_chain[391]));
    BUFFD20BWP7T30P140 delay_inst392 (.I(delay_chain[391]), .Z(delay_chain[392]));
    BUFFD20BWP7T30P140 delay_inst393 (.I(delay_chain[392]), .Z(delay_chain[393]));
    BUFFD20BWP7T30P140 delay_inst394 (.I(delay_chain[393]), .Z(delay_chain[394]));
    BUFFD20BWP7T30P140 delay_inst395 (.I(delay_chain[394]), .Z(delay_chain[395]));
    BUFFD20BWP7T30P140 delay_inst396 (.I(delay_chain[395]), .Z(delay_chain[396]));
    BUFFD20BWP7T30P140 delay_inst397 (.I(delay_chain[396]), .Z(delay_chain[397]));
    BUFFD20BWP7T30P140 delay_inst398 (.I(delay_chain[397]), .Z(delay_chain[398]));
    BUFFD20BWP7T30P140 delay_inst399 (.I(delay_chain[398]), .Z(delay_chain[399]));
    BUFFD20BWP7T30P140 delay_inst400 (.I(delay_chain[399]), .Z(delay_chain[400]));
    BUFFD20BWP7T30P140 delay_inst401 (.I(delay_chain[400]), .Z(delay_chain[401]));
    BUFFD20BWP7T30P140 delay_inst402 (.I(delay_chain[401]), .Z(delay_chain[402]));
    BUFFD20BWP7T30P140 delay_inst403 (.I(delay_chain[402]), .Z(delay_chain[403]));
    BUFFD20BWP7T30P140 delay_inst404 (.I(delay_chain[403]), .Z(delay_chain[404]));
    BUFFD20BWP7T30P140 delay_inst405 (.I(delay_chain[404]), .Z(delay_chain[405]));
    BUFFD20BWP7T30P140 delay_inst406 (.I(delay_chain[405]), .Z(delay_chain[406]));
    BUFFD20BWP7T30P140 delay_inst407 (.I(delay_chain[406]), .Z(delay_chain[407]));
    BUFFD20BWP7T30P140 delay_inst408 (.I(delay_chain[407]), .Z(delay_chain[408]));
    BUFFD20BWP7T30P140 delay_inst409 (.I(delay_chain[408]), .Z(delay_chain[409]));
    BUFFD20BWP7T30P140 delay_inst410 (.I(delay_chain[409]), .Z(delay_chain[410]));
    BUFFD20BWP7T30P140 delay_inst411 (.I(delay_chain[410]), .Z(delay_chain[411]));
    BUFFD20BWP7T30P140 delay_inst412 (.I(delay_chain[411]), .Z(delay_chain[412]));
    BUFFD20BWP7T30P140 delay_inst413 (.I(delay_chain[412]), .Z(delay_chain[413]));
    BUFFD20BWP7T30P140 delay_inst414 (.I(delay_chain[413]), .Z(delay_chain[414]));
    BUFFD20BWP7T30P140 delay_inst415 (.I(delay_chain[414]), .Z(delay_chain[415]));
    BUFFD20BWP7T30P140 delay_inst416 (.I(delay_chain[415]), .Z(delay_chain[416]));
    BUFFD20BWP7T30P140 delay_inst417 (.I(delay_chain[416]), .Z(delay_chain[417]));
    BUFFD20BWP7T30P140 delay_inst418 (.I(delay_chain[417]), .Z(delay_chain[418]));
    BUFFD20BWP7T30P140 delay_inst419 (.I(delay_chain[418]), .Z(delay_chain[419]));
    BUFFD20BWP7T30P140 delay_inst420 (.I(delay_chain[419]), .Z(delay_chain[420]));
    BUFFD20BWP7T30P140 delay_inst421 (.I(delay_chain[420]), .Z(delay_chain[421]));
    BUFFD20BWP7T30P140 delay_inst422 (.I(delay_chain[421]), .Z(delay_chain[422]));
    BUFFD20BWP7T30P140 delay_inst423 (.I(delay_chain[422]), .Z(delay_chain[423]));
    BUFFD20BWP7T30P140 delay_inst424 (.I(delay_chain[423]), .Z(delay_chain[424]));
    BUFFD20BWP7T30P140 delay_inst425 (.I(delay_chain[424]), .Z(delay_chain[425]));
    BUFFD20BWP7T30P140 delay_inst426 (.I(delay_chain[425]), .Z(delay_chain[426]));
    BUFFD20BWP7T30P140 delay_inst427 (.I(delay_chain[426]), .Z(delay_chain[427]));
    BUFFD20BWP7T30P140 delay_inst428 (.I(delay_chain[427]), .Z(delay_chain[428]));
    BUFFD20BWP7T30P140 delay_inst429 (.I(delay_chain[428]), .Z(delay_chain[429]));
    BUFFD20BWP7T30P140 delay_inst430 (.I(delay_chain[429]), .Z(delay_chain[430]));
    BUFFD20BWP7T30P140 delay_inst431 (.I(delay_chain[430]), .Z(delay_chain[431]));
    BUFFD20BWP7T30P140 delay_inst432 (.I(delay_chain[431]), .Z(delay_chain[432]));
    BUFFD20BWP7T30P140 delay_inst433 (.I(delay_chain[432]), .Z(delay_chain[433]));
    BUFFD20BWP7T30P140 delay_inst434 (.I(delay_chain[433]), .Z(delay_chain[434]));
    BUFFD20BWP7T30P140 delay_inst435 (.I(delay_chain[434]), .Z(delay_chain[435]));
    BUFFD20BWP7T30P140 delay_inst436 (.I(delay_chain[435]), .Z(delay_chain[436]));
    BUFFD20BWP7T30P140 delay_inst437 (.I(delay_chain[436]), .Z(delay_chain[437]));
    BUFFD20BWP7T30P140 delay_inst438 (.I(delay_chain[437]), .Z(delay_chain[438]));
    BUFFD20BWP7T30P140 delay_inst439 (.I(delay_chain[438]), .Z(delay_chain[439]));
    BUFFD20BWP7T30P140 delay_inst440 (.I(delay_chain[439]), .Z(delay_chain[440]));
    BUFFD20BWP7T30P140 delay_inst441 (.I(delay_chain[440]), .Z(delay_chain[441]));
    BUFFD20BWP7T30P140 delay_inst442 (.I(delay_chain[441]), .Z(delay_chain[442]));
    BUFFD20BWP7T30P140 delay_inst443 (.I(delay_chain[442]), .Z(delay_chain[443]));
    BUFFD20BWP7T30P140 delay_inst444 (.I(delay_chain[443]), .Z(delay_chain[444]));
    BUFFD20BWP7T30P140 delay_inst445 (.I(delay_chain[444]), .Z(delay_chain[445]));
    BUFFD20BWP7T30P140 delay_inst446 (.I(delay_chain[445]), .Z(delay_chain[446]));
    BUFFD20BWP7T30P140 delay_inst447 (.I(delay_chain[446]), .Z(delay_chain[447]));
    BUFFD20BWP7T30P140 delay_inst448 (.I(delay_chain[447]), .Z(delay_chain[448]));
    BUFFD20BWP7T30P140 delay_inst449 (.I(delay_chain[448]), .Z(delay_chain[449]));
    BUFFD20BWP7T30P140 delay_inst450 (.I(delay_chain[449]), .Z(delay_chain[450]));
    BUFFD20BWP7T30P140 delay_inst451 (.I(delay_chain[450]), .Z(delay_chain[451]));
    BUFFD20BWP7T30P140 delay_inst452 (.I(delay_chain[451]), .Z(delay_chain[452]));
    BUFFD20BWP7T30P140 delay_inst453 (.I(delay_chain[452]), .Z(delay_chain[453]));
    BUFFD20BWP7T30P140 delay_inst454 (.I(delay_chain[453]), .Z(delay_chain[454]));
    BUFFD20BWP7T30P140 delay_inst455 (.I(delay_chain[454]), .Z(delay_chain[455]));
    BUFFD20BWP7T30P140 delay_inst456 (.I(delay_chain[455]), .Z(delay_chain[456]));
    BUFFD20BWP7T30P140 delay_inst457 (.I(delay_chain[456]), .Z(delay_chain[457]));
    BUFFD20BWP7T30P140 delay_inst458 (.I(delay_chain[457]), .Z(delay_chain[458]));
    BUFFD20BWP7T30P140 delay_inst459 (.I(delay_chain[458]), .Z(delay_chain[459]));
    BUFFD20BWP7T30P140 delay_inst460 (.I(delay_chain[459]), .Z(delay_chain[460]));
    BUFFD20BWP7T30P140 delay_inst461 (.I(delay_chain[460]), .Z(delay_chain[461]));
    BUFFD20BWP7T30P140 delay_inst462 (.I(delay_chain[461]), .Z(delay_chain[462]));
    BUFFD20BWP7T30P140 delay_inst463 (.I(delay_chain[462]), .Z(delay_chain[463]));
    BUFFD20BWP7T30P140 delay_inst464 (.I(delay_chain[463]), .Z(delay_chain[464]));
    BUFFD20BWP7T30P140 delay_inst465 (.I(delay_chain[464]), .Z(delay_chain[465]));
    BUFFD20BWP7T30P140 delay_inst466 (.I(delay_chain[465]), .Z(delay_chain[466]));
    BUFFD20BWP7T30P140 delay_inst467 (.I(delay_chain[466]), .Z(delay_chain[467]));
    BUFFD20BWP7T30P140 delay_inst468 (.I(delay_chain[467]), .Z(delay_chain[468]));
    BUFFD20BWP7T30P140 delay_inst469 (.I(delay_chain[468]), .Z(delay_chain[469]));
    BUFFD20BWP7T30P140 delay_inst470 (.I(delay_chain[469]), .Z(delay_chain[470]));
    BUFFD20BWP7T30P140 delay_inst471 (.I(delay_chain[470]), .Z(delay_chain[471]));
    BUFFD20BWP7T30P140 delay_inst472 (.I(delay_chain[471]), .Z(delay_chain[472]));
    BUFFD20BWP7T30P140 delay_inst473 (.I(delay_chain[472]), .Z(delay_chain[473]));
    BUFFD20BWP7T30P140 delay_inst474 (.I(delay_chain[473]), .Z(delay_chain[474]));
    BUFFD20BWP7T30P140 delay_inst475 (.I(delay_chain[474]), .Z(delay_chain[475]));
    BUFFD20BWP7T30P140 delay_inst476 (.I(delay_chain[475]), .Z(delay_chain[476]));
    BUFFD20BWP7T30P140 delay_inst477 (.I(delay_chain[476]), .Z(delay_chain[477]));
    BUFFD20BWP7T30P140 delay_inst478 (.I(delay_chain[477]), .Z(delay_chain[478]));
    BUFFD20BWP7T30P140 delay_inst479 (.I(delay_chain[478]), .Z(delay_chain[479]));
    BUFFD20BWP7T30P140 delay_inst480 (.I(delay_chain[479]), .Z(delay_chain[480]));
    BUFFD20BWP7T30P140 delay_inst481 (.I(delay_chain[480]), .Z(delay_chain[481]));
    BUFFD20BWP7T30P140 delay_inst482 (.I(delay_chain[481]), .Z(delay_chain[482]));
    BUFFD20BWP7T30P140 delay_inst483 (.I(delay_chain[482]), .Z(delay_chain[483]));
    BUFFD20BWP7T30P140 delay_inst484 (.I(delay_chain[483]), .Z(delay_chain[484]));
    BUFFD20BWP7T30P140 delay_inst485 (.I(delay_chain[484]), .Z(delay_chain[485]));
    BUFFD20BWP7T30P140 delay_inst486 (.I(delay_chain[485]), .Z(delay_chain[486]));
    BUFFD20BWP7T30P140 delay_inst487 (.I(delay_chain[486]), .Z(delay_chain[487]));
    BUFFD20BWP7T30P140 delay_inst488 (.I(delay_chain[487]), .Z(delay_chain[488]));
    BUFFD20BWP7T30P140 delay_inst489 (.I(delay_chain[488]), .Z(delay_chain[489]));
    BUFFD20BWP7T30P140 delay_inst490 (.I(delay_chain[489]), .Z(delay_chain[490]));
    BUFFD20BWP7T30P140 delay_inst491 (.I(delay_chain[490]), .Z(delay_chain[491]));
    BUFFD20BWP7T30P140 delay_inst492 (.I(delay_chain[491]), .Z(delay_chain[492]));
    BUFFD20BWP7T30P140 delay_inst493 (.I(delay_chain[492]), .Z(delay_chain[493]));
    BUFFD20BWP7T30P140 delay_inst494 (.I(delay_chain[493]), .Z(delay_chain[494]));
    BUFFD20BWP7T30P140 delay_inst495 (.I(delay_chain[494]), .Z(delay_chain[495]));
    BUFFD20BWP7T30P140 delay_inst496 (.I(delay_chain[495]), .Z(delay_chain[496]));
    BUFFD20BWP7T30P140 delay_inst497 (.I(delay_chain[496]), .Z(delay_chain[497]));
    BUFFD20BWP7T30P140 delay_inst498 (.I(delay_chain[497]), .Z(delay_chain[498]));
    BUFFD20BWP7T30P140 delay_inst499 (.I(delay_chain[498]), .Z(delay_chain[499]));
    BUFFD20BWP7T30P140 delay_inst500 (.I(delay_chain[499]), .Z(delay_chain[500]));
    BUFFD20BWP7T30P140 delay_inst501 (.I(delay_chain[500]), .Z(delay_chain[501]));
    BUFFD20BWP7T30P140 delay_inst502 (.I(delay_chain[501]), .Z(delay_chain[502]));
    BUFFD20BWP7T30P140 delay_inst503 (.I(delay_chain[502]), .Z(delay_chain[503]));
    BUFFD20BWP7T30P140 delay_inst504 (.I(delay_chain[503]), .Z(delay_chain[504]));
    BUFFD20BWP7T30P140 delay_inst505 (.I(delay_chain[504]), .Z(delay_chain[505]));
    BUFFD20BWP7T30P140 delay_inst506 (.I(delay_chain[505]), .Z(delay_chain[506]));
    BUFFD20BWP7T30P140 delay_inst507 (.I(delay_chain[506]), .Z(delay_chain[507]));
    BUFFD20BWP7T30P140 delay_inst508 (.I(delay_chain[507]), .Z(delay_chain[508]));
    BUFFD20BWP7T30P140 delay_inst509 (.I(delay_chain[508]), .Z(delay_chain[509]));
    BUFFD20BWP7T30P140 delay_inst510 (.I(delay_chain[509]), .Z(delay_chain[510]));
    BUFFD20BWP7T30P140 delay_inst511 (.I(delay_chain[510]), .Z(delay_chain[511]));
endmodule
